LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Or2 IS
  PORT (
    X, Y : IN  STD_ULOGIC;
    Z    : OUT STD_ULOGIC
  );
END ENTITY Or2;

ARCHITECTURE ImplOr2 OF Or2 IS
  BEGIN
    Z <= X OR Y;
END ARCHITECTURE ImplOr2;
